module connect4(

);